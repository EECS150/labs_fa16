module full_adder (
    input a,
    input b,
    input carry_in,
    output sum, 
    output carry_out
);

    // Insert your RTL here to calculate the sum and carry out bits
    
    // Remove these assign statements once you write your own RTL
    assign sum = 1'b0;
    assign carry_out = 1'b0;

endmodule