module tone_generator (
    input output_enable,
    input [23:0] tone_switch_period, 
    input clk,
    input rst,
    output square_wave_out
);

    // Remove this line once you have copied over your tone_generator implementation
    assign square_wave_out = 0;

endmodule
