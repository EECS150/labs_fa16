module structural_adder (
    input [3:0] a,
    input [3:0] b,
    output [4:0] sum
);

    // Instantiate your full adder cells here and wire them together

    // Remove this line when you've added your own RTL
    assign sum = 5'b0;
endmodule