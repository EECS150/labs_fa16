module music_streamer (
    input clk,
    input [1:0] tempo,
    input pause,
    output [23:0] tone
);

endmodule
